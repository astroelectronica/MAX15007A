.title KiCad schematic
.include "C:/AE/MAX15007A/_models/C2012X7R2A104K125AA_p.mod"
.include "C:/AE/MAX15007A/_models/C3216X5R1C106M160AA_p.mod"
.include "C:/AE/MAX15007A/_models/C3216X7R2A105M160AA_p.mod"
.include "C:/AE/MAX15007A/_models/MAX15007A.lib"
V1 /VIN 0 {VSOURCE}
XU3 /VIN 0 C2012X7R2A104K125AA_p
R1 /VIN /EN {REN}
XU2 /VIN 0 C3216X7R2A105M160AA_p
I1 /VOUT 0 {ILOAD}
XU5 /VOUT 0 C2012X7R2A104K125AA_p
XU4 /VOUT 0 C3216X5R1C106M160AA_p
XU1 /VIN unconnected-_U1-NC-Pad2_ /EN unconnected-_U1-NC-Pad4_ 0 unconnected-_U1-NC-Pad6_ unconnected-_U1-NC-Pad7_ /VOUT MAX15007A
.end
